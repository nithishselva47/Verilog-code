//nithish selva M 20l136//
module halfadder(
    input a,b,
    output s,co
    );
assign s=a^b;
  assign co=a&b;
endmodule
